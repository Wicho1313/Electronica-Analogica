** Profile: "SCHEMATIC1-MediaOnda_Filtro"  [ C:\Users\Wicho\Documents\ESCOM\Analogica\Practicas\P02\MediaOnda_Filtro-PSpiceFiles\SCHEMATIC1\MediaOnda_Filtro.sim ] 

** Creating circuit file "MediaOnda_Filtro.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Wicho\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 60ms 0 50u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
